module seven_seg_decodera(F, I);
	input [3:0] I;
	output [6:0] F;
	
	reg [6:0] F;
	
	always @(I) begin
		case ({I})
			4'b0000: F = 7'b0000001;
			4'b0001: F = 7'b1001111;
			4'b0010: F = 7'b0010010;
			4'b0011: F = 7'b0000110;
			4'b0100: F = 7'b1001100;
			4'b0101: F = 7'b0100100;
			4'b0110: F = 7'b0100000;
			4'b0111: F = 7'b0001111;
			4'b1000: F = 7'b0000000;
			4'b1001: F = 7'b0000100;
			4'b1010: F = 7'b0001000;
			4'b1011: F = 7'b1100000;
			4'b1100: F = 7'b0110001;
			4'b1101: F = 7'b1000010;
			4'b1110: F = 7'b0110000;
			4'b1111: F = 7'b0111000;
		endcase
	end
endmodule
	